module main

struct Note {
	text string
}
