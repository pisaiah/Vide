module main

import iui as ui
import gg
