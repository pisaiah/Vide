// Console Hider - Public Domain
module hc

pub fn hide_console_win() {
}
